//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/01/2018 07:47:04 PM
// Design Name: 
// Module Name: crosswalk
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module crosswalk(
    output reg walk_light,
    output reg stop_light,
    input red_trffc_light,
    input ylw_trffc_light,
    input clk    
);
endmodule
